`define CONFIG_DIFFTEST_INTERFACE_WIDTH 33363
`define CONFIG_DIFFTEST_STEPWIDTH 7
`define CONFIG_DIFFTEST_BATCH_IO_WITDH 16000
`define CONFIG_DIFFTEST_DEFERRED_RESULT
`define CONFIG_DIFFTEST_INTERNAL_STEP
`define CONFIG_DIFFTEST_FPGA
`define CONFIG_DIFFTEST_CLOCKGATE
`define CPU_XIANGSHAN
