
module array_0_2_ext(
  input RW0_clk,
  input [12:0] RW0_addr,
  input RW0_en,
  input RW0_wmode,
  input [4:0] RW0_wdata,
  output [4:0] RW0_rdata
);

  reg reg_RW0_ren;
  reg [12:0] reg_RW0_addr;
  (* ram_style = "ultra" *) reg [4:0] ram [8191:0];
  `ifdef RANDOMIZE_MEM_INIT
    integer initvar;
    initial begin
      #`RANDOMIZE_DELAY begin end
      for (initvar = 0; initvar < 8192; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
      reg_RW0_addr = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge RW0_clk)
    reg_RW0_ren <= RW0_en && !RW0_wmode;
  always @(posedge RW0_clk)
    if (RW0_en && !RW0_wmode) reg_RW0_addr <= RW0_addr;
  always @(posedge RW0_clk)
    if (RW0_en && RW0_wmode) begin
      for (i=0;i<1;i=i+1) begin
        ram[RW0_addr][i*5 +: 5] <= RW0_wdata[i*5 +: 5];
      end
    end
  `ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] RW0_random;
  `ifdef RANDOMIZE_MEM_INIT
    initial begin
      #`RANDOMIZE_DELAY begin end
      RW0_random = {$random};
      reg_RW0_ren = RW0_random[0];
    end
  `endif
  always @(posedge RW0_clk) RW0_random <= {$random};
  assign RW0_rdata = reg_RW0_ren ? ram[reg_RW0_addr] : RW0_random[4:0];
  `else
  assign RW0_rdata = ram[reg_RW0_addr];
  `endif

endmodule